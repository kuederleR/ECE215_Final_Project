module FrequencyDetector();

endmodule
